module Top (
	input i_rst_n,
	input i_clk,
	// choose different states 
	input i_key_0,   // reset
	input i_key_1,	 // start or stop
	input i_key_2,	 // play and pause
	
	// OUR SWITCHES 
	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************
	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************
	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************
	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************
	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************


	input i_play_or_record, // switch SW[0] 0 for record 1 for playing

	input i_speed_control, // switch SW[1]  1 for fast, 0 for slow

	input i_speed_b0, // switch SW[2-4]  choose up/down sample rate 1-8
	input i_speed_b1,
	input i_speed_b2,
	input i_order,


	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************
	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************
	//  REMEMBER TO CHANGE DE2_115 *******************************************************************************
	output [2:0] o_top_state,
	output o_LEDG,
	output [3:0] o_LEDR,
	output [3:0] o_record_LED,
	output [3:0] o_play_LED,
	output [5:0] o_time,
	// input [3:0] i_speed, // design how user can decide mode on your own
	
	// AudDSP and SRAM
	output [19:0] o_SRAM_ADDR,
	inout  [15:0] io_SRAM_DQ,
	output        o_SRAM_WE_N, // **** enable ****
	output        o_SRAM_CE_N, // dont care about these 
	output        o_SRAM_OE_N, //
 	output        o_SRAM_LB_N, //
	output        o_SRAM_UB_N, // all default settings
	
	// I2C
	input  i_clk_100k, 
	output o_I2C_SCLK,
	inout  io_I2C_SDAT,
	
	// AudPlayer
	inout  i_AUD_BCLK,

	input  i_AUD_ADCDAT,    // FROM RECORDER: analog to digital -> store inside sram
	inout  i_AUD_ADCLRCK,	// recieving from WM8731

	
	inout  i_AUD_DACLRCK,	// FOR PLAYER: digital to analog -> 
	output o_AUD_DACDAT		// outputting to WM8731

	// SEVENDECODER (optional display)
	// output [5:0] o_record_time,
	// output [5:0] o_play_time,

	// LCD (optional display)
	// input        i_clk_800k,
	// inout  [7:0] o_LCD_DATA,
	// output       o_LCD_EN,
	// output       o_LCD_RS,
	// output       o_LCD_RW,
	// output       o_LCD_ON,
	// output       o_LCD_BLON,

	// LED
	// output  [8:0] o_ledg,
	// output [17:0] o_ledr
);

// design the FSM and states as you like
parameter S_IDLE       = 0;
parameter S_I2C        = 1;
parameter S_RECD       = 2;
//parameter S_RECD_PAUSE = 3;
parameter S_PLAY       = 3;
parameter S_PLAY_PAUSE = 4;

logic i2c_oen, i2c_sdat;
logic [19:0] addr_record, addr_play;
logic [15:0] data_record, data_play, dac_data;
logic ledg_r, ledg_w;
logic [3:0] ledr_r, ledr_w;
logic [3:0] led_record;
logic [3:0] led_play;
logic [2:0] five_dec_r, five_dec_w;

// below is a simple example for module division
// you can design these as you like


// register decleration
logic [2:0] state_w, state_r;
logic I2C_start_w, I2C_start_r; 
logic PLAYER_start_w, PLAYER_start_r;
logic RECORDER_start_w, RECORDER_start_r;
logic [5:0] run_time_r;
logic [5:0] play_time;
// wire delcaration
wire I2C_done, play_done, record_done;
// === I2cInitializer ===
// sequentially sent out settings to initialize WM8731 with I2C protocal
I2cInitializer init0(
	.i_rst_n(i_rst_n),
	.i_clk(i_clk_100k),
	.i_start(I2C_start_r),
	.o_finished(I2C_done),
	.o_sclk(o_I2C_SCLK),
	.o_sdat(io_I2C_SDAT),
	.o_oen(i2c_oen) // you are outputing (you are not outputing only when you are "ack"ing.)
);

// === AudDSP ===
// responsible for DSP operations including fast play and slow play at different speed
// in other words, determine which data addr to be fetch for player 
// AudDSP dsp0(
// 	.i_rst_n(i_rst_n),
// 	.i_clk(i_clk),
// 	.i_start(),
// 	.i_pause(),
// 	.i_stop(),
// 	.i_speed(),
// 	.i_fast(),
// 	.i_slow_0(), // constant interpolation
// 	.i_slow_1(), // linear interpolation
// 	.i_daclrck(i_AUD_DACLRCK),
// 	.i_sram_data(data_play),
// 	.o_dac_data(dac_data),
// 	.o_sram_addr(addr_play)
// );

// === AudPlayer ===
// receive data address from DSP and fetch data to sent to WM8731 with I2S protocal
AudPlayer player0(
	.i_rst_n(i_rst_n),
	.i_bclk(i_AUD_BCLK),
	.i_daclrck(i_AUD_DACLRCK), // left right channel
	.i_speed({i_speed_control, i_speed_b2, i_speed_b1, i_speed_b0}), // playback speed
	.i_start(PLAYER_start_r), //start or stop
	.i_pause(i_key_2), // play or pause
	// .i_en(), // enable AudPlayer only when playing audio, work with AudDSP
	.i_dac_data(data_play), //dac_data from sram
	.o_aud_dacdat(o_AUD_DACDAT), //result for WM8731
	//.o_aud_dacdat(player_out),
	.o_sram_addr(addr_play), //addr player want from sram
	.o_done(play_done),
	.o_led(led_play),
	.o_play_time(play_time),
	.i_order(i_order)
);

// === AudRecorder ===
// receive data from WM8731 with I2S protocal and save to SRAM
AudRecorder recorder0(
	.i_rst_n(i_rst_n), 
	.i_clk(i_AUD_BCLK),
	.i_lrc(i_AUD_ADCLRCK), // left/right channel
	.i_start(RECORDER_start_r), // once it start, record 32 sec
	.i_data(i_AUD_ADCDAT), // data from WM8731
	.o_address(addr_record), // addr to sram
	.o_data(data_record), //data to sram
	.o_run_time(run_time_r),
	// OUR CONTROLS
	.o_done(record_done),
	.o_led(led_record),
	.o_SRAM_WE(o_SRAM_WE_N)
);


// Recorder adc(
// 	.i_rst_n(i_rst_n), 
// 	.i_record(RECORDER_start_r), 
// 	.i_ADCLRCK(i_AUD_ADCLRCK), 
// 	.i_ADCDAT(i_AUD_ADCDAT), 
// 	.i_BCLK(i_AUD_BCLK), 
// 	.o_SRAM_WE(o_SRAM_WE_N),
// 	.o_SRAM_DATA(data_record), 
// 	.o_done(record_done), 
// 	.SRAM_ADDR(addr_record), 
// 	.o_REC_STATE()
// );

// === FINITE　STATE MACHINE ===
always_comb begin
	state_w = state_r;
	ledr_w = ledr_r;
	ledg_w = 1;
	five_dec_w = five_dec_r;
	case (state_r)
		S_I2C: begin
			ledr_w = 4'b0000;
			// start I2C
			// 1. I2C start on
			// 2. Wait for I2C done signal
			// 3. Go to S_IDLE
			if(I2C_done)begin
				state_w = S_IDLE;
			end

		end
		S_IDLE: begin
			five_dec_w = 3'd0;
			ledr_w = 1;
			// wait for record / play control switch (key 1)
			// if record -> next state = S_RECD
			// if play -> next state = S_PLAY
			// else -> stay in S_IDLE
			if(i_key_1)begin // start
				if (i_play_or_record) begin
					state_w = S_PLAY;
				end else begin
					state_w = S_RECD;
				end
			end
		end
		
		S_RECD: begin
			ledr_w = 4'b0010;
			five_dec_w = 3'd2;
			//If finish recording go back to S_IDLE
			if (record_done) begin
				state_w = S_IDLE;
			end

		end
		S_PLAY: begin
			ledr_w = 4'b011;
			five_dec_w = 3'd1;
			// If finish playing go back to S_IDLE
			// If pause then go to S_PLAY_PAUSE
			if (play_done) begin // finish
				state_w = S_IDLE;
			end else if (i_key_2) begin //pause
				state_w = S_PLAY_PAUSE;
			end else if (i_key_1) begin // stop
				state_w = S_IDLE;
			end else begin
				state_w = S_PLAY;
			end
		end
		S_PLAY_PAUSE: begin
			ledr_w = 4'd4;
			five_dec_w = 3'd3;
			if(i_key_2)begin
				state_w = S_PLAY;
			end
			
		end
		default: begin
			ledr_w = 4'b1111;
			ledg_w = 1;
		end
	endcase
	if (i_key_0) begin
		state_w = S_I2C;
	end
end



always_comb begin
	// design your control here
	RECORDER_start_w = RECORDER_start_r;
	PLAYER_start_w = PLAYER_start_r;
	I2C_start_w = I2C_start_r;
	case (state_r)
		S_I2C: begin
			I2C_start_w = 1;
			if (I2C_done) begin
				I2C_start_w = 0;
			end
		end
		S_IDLE: begin
			I2C_start_w = 0;
			RECORDER_start_w = 0;
			PLAYER_start_w = 0;
		end
		S_RECD: begin
			PLAYER_start_w = 0;
			RECORDER_start_w = 1;
		end
		S_PLAY: begin
			PLAYER_start_w = 1;
			RECORDER_start_w = 0;
		end
		S_PLAY_PAUSE: begin
		end
		default: begin
			
		end
	endcase
	// if (i_key_0) begin
	// 	PLAYER_start_w = 0;
	// 	RECORDER_start_w = 0;
	// end
end

always_ff @(posedge i_clk or negedge i_rst_n) begin
	if (!i_rst_n) begin
		RECORDER_start_r <=0;
		PLAYER_start_r <=0;
		state_r <= S_I2C;
		I2C_start_r <= 1;
		ledr_r <=4'b1000;
		ledg_r <=1;
		five_dec_r <=0;
		// run_time_r <= 0;
	end
	else begin
		RECORDER_start_r <=RECORDER_start_w;
		PLAYER_start_r <= PLAYER_start_w;
		state_r <= state_w;
		I2C_start_r <=  I2C_start_w;
		ledg_r <= ledg_w;
		ledr_r <= ledr_w;
		five_dec_r <=five_dec_w;
		// run_time_r <= run_time_w;
	end
end
//assign io_I2C_SDAT = (i2c_oen) ? i2c_sdat : 1'bz;

assign o_SRAM_ADDR = (state_r == S_PLAY) ? addr_play[19:0] : addr_record ;
assign io_SRAM_DQ  = (state_r == S_PLAY) ?  16'dz : data_record; // sram_dq as output
assign data_play   = (state_r == S_PLAY) ? io_SRAM_DQ : 16'dz; // sram_dq as input
assign o_time      = (state_r == S_RECD) ? run_time_r : ((state_r == S_PLAY || state_r == S_PLAY_PAUSE) ? play_time : 0);
//assign o_SRAM_WE_N = (state_r == S_RECD) ? 1'b0 : 1'b1; // if recording than set 0 to write data, else set 1 to read
assign o_SRAM_CE_N = 1'b0;
assign o_SRAM_OE_N = 1'b0;
assign o_SRAM_LB_N = 1'b0;
assign o_SRAM_UB_N = 1'b0;
assign o_LEDR = ledr_r;
assign o_LEDG = ledg_r;
assign o_record_LED = led_record;
assign o_play_LED = led_play;
assign o_top_state = five_dec_r;

// assign o_AUD_DACDAT = (player_state == ) ? player_out : 1'bz;
endmodule

