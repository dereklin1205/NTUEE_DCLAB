task change_view;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[1];
  o_c_state[1] = i_c_state[2];
  o_c_state[2] = i_c_state[3];
  o_c_state[3] = i_c_state[0];
  o_c_state[4] = i_c_state[22];
  o_c_state[5] = i_c_state[11];
  o_c_state[6] = i_c_state[7];
  o_c_state[7] = i_c_state[8];
  o_c_state[8] = i_c_state[9];
  o_c_state[9] = i_c_state[6];
  o_c_state[10] = i_c_state[4];
  o_c_state[11] = i_c_state[17];
  o_c_state[12] = i_c_state[13];
  o_c_state[13] = i_c_state[14];
  o_c_state[14] = i_c_state[15];
  o_c_state[15] = i_c_state[12];
  o_c_state[16] = i_c_state[10];
  o_c_state[17] = i_c_state[23];
  o_c_state[18] = i_c_state[19];
  o_c_state[19] = i_c_state[20];
  o_c_state[20] = i_c_state[21];
  o_c_state[21] = i_c_state[18];
  o_c_state[22] = i_c_state[16];
  o_c_state[23] = i_c_state[5];
  o_c_state[24] = i_c_state[25];
  o_c_state[25] = i_c_state[26];
  o_c_state[26] = i_c_state[27];
  o_c_state[27] = i_c_state[24];
  o_c_state[28] = i_c_state[46];
  o_c_state[29] = i_c_state[35];
  o_c_state[30] = i_c_state[31];
  o_c_state[31] = i_c_state[32];
  o_c_state[32] = i_c_state[33];
  o_c_state[33] = i_c_state[30];
  o_c_state[34] = i_c_state[28];
  o_c_state[35] = i_c_state[41];
  o_c_state[36] = i_c_state[37];
  o_c_state[37] = i_c_state[38];
  o_c_state[38] = i_c_state[39];
  o_c_state[39] = i_c_state[36];
  o_c_state[40] = i_c_state[34];
  o_c_state[41] = i_c_state[47];
  o_c_state[42] = i_c_state[43];
  o_c_state[43] = i_c_state[44];
  o_c_state[44] = i_c_state[45];
  o_c_state[45] = i_c_state[42];
  o_c_state[46] = i_c_state[40];
  o_c_state[47] = i_c_state[29];
  end
  endtask
task Front_clockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[6] = i_c_state[0];
  o_c_state[11] = i_c_state[1];
  o_c_state[2] = i_c_state[2];
  o_c_state[3] = i_c_state[3];
  o_c_state[4] = i_c_state[4];
  o_c_state[9] = i_c_state[5];
  o_c_state[12] = i_c_state[6];
  o_c_state[7] = i_c_state[7];
  o_c_state[8] = i_c_state[8];
  o_c_state[16] = i_c_state[9];
  o_c_state[10] = i_c_state[10];
  o_c_state[15] = i_c_state[11];
  o_c_state[18] = i_c_state[12];
  o_c_state[13] = i_c_state[13];
  o_c_state[14] = i_c_state[14];
  o_c_state[22] = i_c_state[15];
  o_c_state[19] = i_c_state[16];
  o_c_state[17] = i_c_state[17];
  o_c_state[0] = i_c_state[18];
  o_c_state[5] = i_c_state[19];
  o_c_state[20] = i_c_state[20];
  o_c_state[21] = i_c_state[21];
  o_c_state[1] = i_c_state[22];
  o_c_state[23] = i_c_state[23];
  o_c_state[30] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[28];
  o_c_state[33] = i_c_state[29];
  o_c_state[36] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[40] = i_c_state[33];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[42] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[39];
  o_c_state[43] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[24] = i_c_state[42];
  o_c_state[29] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Front_counterclockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[18] = i_c_state[0];
  o_c_state[22] = i_c_state[1];
  o_c_state[2] = i_c_state[2];
  o_c_state[3] = i_c_state[3];
  o_c_state[4] = i_c_state[4];
  o_c_state[19] = i_c_state[5];
  o_c_state[0] = i_c_state[6];
  o_c_state[7] = i_c_state[7];
  o_c_state[8] = i_c_state[8];
  o_c_state[5] = i_c_state[9];
  o_c_state[10] = i_c_state[10];
  o_c_state[1] = i_c_state[11];
  o_c_state[6] = i_c_state[12];
  o_c_state[13] = i_c_state[13];
  o_c_state[14] = i_c_state[14];
  o_c_state[11] = i_c_state[15];
  o_c_state[9] = i_c_state[16];
  o_c_state[17] = i_c_state[17];
  o_c_state[12] = i_c_state[18];
  o_c_state[16] = i_c_state[19];
  o_c_state[20] = i_c_state[20];
  o_c_state[21] = i_c_state[21];
  o_c_state[15] = i_c_state[22];
  o_c_state[23] = i_c_state[23];
  o_c_state[42] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[28];
  o_c_state[43] = i_c_state[29];
  o_c_state[24] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[29] = i_c_state[33];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[30] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[39];
  o_c_state[33] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[36] = i_c_state[42];
  o_c_state[40] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Left_clockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[4];
  o_c_state[1] = i_c_state[1];
  o_c_state[2] = i_c_state[2];
  o_c_state[3] = i_c_state[21];
  o_c_state[4] = i_c_state[14];
  o_c_state[5] = i_c_state[0];
  o_c_state[6] = i_c_state[6];
  o_c_state[7] = i_c_state[7];
  o_c_state[8] = i_c_state[23];
  o_c_state[9] = i_c_state[3];
  o_c_state[10] = i_c_state[10];
  o_c_state[11] = i_c_state[11];
  o_c_state[12] = i_c_state[12];
  o_c_state[13] = i_c_state[13];
  o_c_state[14] = i_c_state[5];
  o_c_state[15] = i_c_state[9];
  o_c_state[16] = i_c_state[16];
  o_c_state[17] = i_c_state[17];
  o_c_state[18] = i_c_state[22];
  o_c_state[19] = i_c_state[19];
  o_c_state[20] = i_c_state[20];
  o_c_state[21] = i_c_state[15];
  o_c_state[22] = i_c_state[8];
  o_c_state[23] = i_c_state[18];
  o_c_state[24] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[45];
  o_c_state[28] = i_c_state[28];
  o_c_state[29] = i_c_state[29];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[47];
  o_c_state[33] = i_c_state[27];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[33];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[42] = i_c_state[46];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[39];
  o_c_state[46] = i_c_state[32];
  o_c_state[47] = i_c_state[42];
  end
  endtask
task Left_counterclockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[5];
  o_c_state[1] = i_c_state[1];
  o_c_state[2] = i_c_state[2];
  o_c_state[3] = i_c_state[9];
  o_c_state[4] = i_c_state[0];
  o_c_state[5] = i_c_state[14];
  o_c_state[6] = i_c_state[6];
  o_c_state[7] = i_c_state[7];
  o_c_state[8] = i_c_state[22];
  o_c_state[9] = i_c_state[15];
  o_c_state[10] = i_c_state[10];
  o_c_state[11] = i_c_state[11];
  o_c_state[12] = i_c_state[12];
  o_c_state[13] = i_c_state[13];
  o_c_state[14] = i_c_state[4];
  o_c_state[15] = i_c_state[21];
  o_c_state[16] = i_c_state[16];
  o_c_state[17] = i_c_state[17];
  o_c_state[18] = i_c_state[23];
  o_c_state[19] = i_c_state[19];
  o_c_state[20] = i_c_state[20];
  o_c_state[21] = i_c_state[3];
  o_c_state[22] = i_c_state[18];
  o_c_state[23] = i_c_state[8];
  o_c_state[24] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[33];
  o_c_state[28] = i_c_state[28];
  o_c_state[29] = i_c_state[29];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[46];
  o_c_state[33] = i_c_state[39];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[45];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[42] = i_c_state[47];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[27];
  o_c_state[46] = i_c_state[42];
  o_c_state[47] = i_c_state[32];
  end
  endtask
task Right_clockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[0];
  o_c_state[7] = i_c_state[1];
  o_c_state[17] = i_c_state[2];
  o_c_state[3] = i_c_state[3];
  o_c_state[4] = i_c_state[4];
  o_c_state[5] = i_c_state[5];
  o_c_state[10] = i_c_state[6];
  o_c_state[13] = i_c_state[7];
  o_c_state[8] = i_c_state[8];
  o_c_state[9] = i_c_state[9];
  o_c_state[20] = i_c_state[10];
  o_c_state[6] = i_c_state[11];
  o_c_state[16] = i_c_state[12];
  o_c_state[19] = i_c_state[13];
  o_c_state[14] = i_c_state[14];
  o_c_state[15] = i_c_state[15];
  o_c_state[2] = i_c_state[16];
  o_c_state[12] = i_c_state[17];
  o_c_state[18] = i_c_state[18];
  o_c_state[1] = i_c_state[19];
  o_c_state[11] = i_c_state[20];
  o_c_state[21] = i_c_state[21];
  o_c_state[22] = i_c_state[22];
  o_c_state[23] = i_c_state[23];
  o_c_state[24] = i_c_state[24];
  o_c_state[31] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[28];
  o_c_state[29] = i_c_state[29];
  o_c_state[34] = i_c_state[30];
  o_c_state[37] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[33] = i_c_state[33];
  o_c_state[44] = i_c_state[34];
  o_c_state[30] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[43] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[39];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[42] = i_c_state[42];
  o_c_state[25] = i_c_state[43];
  o_c_state[35] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Right_counterclockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[0];
  o_c_state[19] = i_c_state[1];
  o_c_state[16] = i_c_state[2];
  o_c_state[3] = i_c_state[3];
  o_c_state[4] = i_c_state[4];
  o_c_state[5] = i_c_state[5];
  o_c_state[11] = i_c_state[6];
  o_c_state[1] = i_c_state[7];
  o_c_state[8] = i_c_state[8];
  o_c_state[9] = i_c_state[9];
  o_c_state[6] = i_c_state[10];
  o_c_state[20] = i_c_state[11];
  o_c_state[17] = i_c_state[12];
  o_c_state[7] = i_c_state[13];
  o_c_state[14] = i_c_state[14];
  o_c_state[15] = i_c_state[15];
  o_c_state[12] = i_c_state[16];
  o_c_state[2] = i_c_state[17];
  o_c_state[18] = i_c_state[18];
  o_c_state[13] = i_c_state[19];
  o_c_state[10] = i_c_state[20];
  o_c_state[21] = i_c_state[21];
  o_c_state[22] = i_c_state[22];
  o_c_state[23] = i_c_state[23];
  o_c_state[24] = i_c_state[24];
  o_c_state[43] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[28];
  o_c_state[29] = i_c_state[29];
  o_c_state[35] = i_c_state[30];
  o_c_state[25] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[33] = i_c_state[33];
  o_c_state[30] = i_c_state[34];
  o_c_state[44] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[31] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[39];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[42] = i_c_state[42];
  o_c_state[37] = i_c_state[43];
  o_c_state[34] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Top_clockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[3] = i_c_state[0];
  o_c_state[0] = i_c_state[1];
  o_c_state[1] = i_c_state[2];
  o_c_state[2] = i_c_state[3];
  o_c_state[10] = i_c_state[4];
  o_c_state[5] = i_c_state[5];
  o_c_state[9] = i_c_state[6];
  o_c_state[6] = i_c_state[7];
  o_c_state[7] = i_c_state[8];
  o_c_state[8] = i_c_state[9];
  o_c_state[16] = i_c_state[10];
  o_c_state[11] = i_c_state[11];
  o_c_state[12] = i_c_state[12];
  o_c_state[13] = i_c_state[13];
  o_c_state[14] = i_c_state[14];
  o_c_state[15] = i_c_state[15];
  o_c_state[22] = i_c_state[16];
  o_c_state[17] = i_c_state[17];
  o_c_state[18] = i_c_state[18];
  o_c_state[19] = i_c_state[19];
  o_c_state[20] = i_c_state[20];
  o_c_state[21] = i_c_state[21];
  o_c_state[4] = i_c_state[22];
  o_c_state[23] = i_c_state[23];
  o_c_state[27] = i_c_state[24];
  o_c_state[24] = i_c_state[25];
  o_c_state[25] = i_c_state[26];
  o_c_state[26] = i_c_state[27];
  o_c_state[34] = i_c_state[28];
  o_c_state[29] = i_c_state[29];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[33] = i_c_state[33];
  o_c_state[40] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[39];
  o_c_state[46] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[42] = i_c_state[42];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[28] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Top_counterclockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[1] = i_c_state[0];
  o_c_state[2] = i_c_state[1];
  o_c_state[3] = i_c_state[2];
  o_c_state[0] = i_c_state[3];
  o_c_state[22] = i_c_state[4];
  o_c_state[5] = i_c_state[5];
  o_c_state[7] = i_c_state[6];
  o_c_state[8] = i_c_state[7];
  o_c_state[9] = i_c_state[8];
  o_c_state[6] = i_c_state[9];
  o_c_state[4] = i_c_state[10];
  o_c_state[11] = i_c_state[11];
  o_c_state[12] = i_c_state[12];
  o_c_state[13] = i_c_state[13];
  o_c_state[14] = i_c_state[14];
  o_c_state[15] = i_c_state[15];
  o_c_state[10] = i_c_state[16];
  o_c_state[17] = i_c_state[17];
  o_c_state[18] = i_c_state[18];
  o_c_state[19] = i_c_state[19];
  o_c_state[20] = i_c_state[20];
  o_c_state[21] = i_c_state[21];
  o_c_state[16] = i_c_state[22];
  o_c_state[23] = i_c_state[23];
  o_c_state[25] = i_c_state[24];
  o_c_state[26] = i_c_state[25];
  o_c_state[27] = i_c_state[26];
  o_c_state[24] = i_c_state[27];
  o_c_state[46] = i_c_state[28];
  o_c_state[29] = i_c_state[29];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[33] = i_c_state[33];
  o_c_state[28] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[38];
  o_c_state[39] = i_c_state[39];
  o_c_state[34] = i_c_state[40];
  o_c_state[41] = i_c_state[41];
  o_c_state[42] = i_c_state[42];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[40] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Down_clockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[0];
  o_c_state[1] = i_c_state[1];
  o_c_state[2] = i_c_state[2];
  o_c_state[3] = i_c_state[3];
  o_c_state[4] = i_c_state[4];
  o_c_state[5] = i_c_state[23];
  o_c_state[6] = i_c_state[6];
  o_c_state[7] = i_c_state[7];
  o_c_state[8] = i_c_state[8];
  o_c_state[9] = i_c_state[9];
  o_c_state[10] = i_c_state[10];
  o_c_state[11] = i_c_state[5];
  o_c_state[12] = i_c_state[15];
  o_c_state[13] = i_c_state[12];
  o_c_state[14] = i_c_state[13];
  o_c_state[15] = i_c_state[14];
  o_c_state[16] = i_c_state[16];
  o_c_state[17] = i_c_state[11];
  o_c_state[18] = i_c_state[21];
  o_c_state[19] = i_c_state[18];
  o_c_state[20] = i_c_state[19];
  o_c_state[21] = i_c_state[20];
  o_c_state[22] = i_c_state[22];
  o_c_state[23] = i_c_state[17];
  o_c_state[24] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[28];
  o_c_state[29] = i_c_state[47];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[33] = i_c_state[33];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[29];
  o_c_state[36] = i_c_state[39];
  o_c_state[37] = i_c_state[36];
  o_c_state[38] = i_c_state[37];
  o_c_state[39] = i_c_state[38];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[35];
  o_c_state[42] = i_c_state[42];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[41];
  end
  endtask
task Down_counterclockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[0];
  o_c_state[1] = i_c_state[1];
  o_c_state[2] = i_c_state[2];
  o_c_state[3] = i_c_state[3];
  o_c_state[4] = i_c_state[4];
  o_c_state[5] = i_c_state[11];
  o_c_state[6] = i_c_state[6];
  o_c_state[7] = i_c_state[7];
  o_c_state[8] = i_c_state[8];
  o_c_state[9] = i_c_state[9];
  o_c_state[10] = i_c_state[10];
  o_c_state[11] = i_c_state[17];
  o_c_state[12] = i_c_state[13];
  o_c_state[13] = i_c_state[14];
  o_c_state[14] = i_c_state[15];
  o_c_state[15] = i_c_state[12];
  o_c_state[16] = i_c_state[16];
  o_c_state[17] = i_c_state[23];
  o_c_state[18] = i_c_state[19];
  o_c_state[19] = i_c_state[20];
  o_c_state[20] = i_c_state[21];
  o_c_state[21] = i_c_state[18];
  o_c_state[22] = i_c_state[22];
  o_c_state[23] = i_c_state[5];
  o_c_state[24] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[26];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[28];
  o_c_state[29] = i_c_state[35];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[31];
  o_c_state[32] = i_c_state[32];
  o_c_state[33] = i_c_state[33];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[41];
  o_c_state[36] = i_c_state[37];
  o_c_state[37] = i_c_state[38];
  o_c_state[38] = i_c_state[39];
  o_c_state[39] = i_c_state[36];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[47];
  o_c_state[42] = i_c_state[42];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[44];
  o_c_state[45] = i_c_state[45];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[29];
  end
  endtask
task Back_clockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[0];
  o_c_state[1] = i_c_state[1];
  o_c_state[2] = i_c_state[20];
  o_c_state[3] = i_c_state[10];
  o_c_state[4] = i_c_state[7];
  o_c_state[5] = i_c_state[5];
  o_c_state[6] = i_c_state[6];
  o_c_state[7] = i_c_state[17];
  o_c_state[8] = i_c_state[2];
  o_c_state[9] = i_c_state[9];
  o_c_state[10] = i_c_state[13];
  o_c_state[11] = i_c_state[11];
  o_c_state[12] = i_c_state[12];
  o_c_state[13] = i_c_state[23];
  o_c_state[14] = i_c_state[8];
  o_c_state[15] = i_c_state[15];
  o_c_state[16] = i_c_state[16];
  o_c_state[17] = i_c_state[21];
  o_c_state[18] = i_c_state[18];
  o_c_state[19] = i_c_state[19];
  o_c_state[20] = i_c_state[14];
  o_c_state[21] = i_c_state[4];
  o_c_state[22] = i_c_state[22];
  o_c_state[23] = i_c_state[3];
  o_c_state[24] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[44];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[31];
  o_c_state[29] = i_c_state[29];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[41];
  o_c_state[32] = i_c_state[26];
  o_c_state[33] = i_c_state[33];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[32];
  o_c_state[39] = i_c_state[39];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[45];
  o_c_state[42] = i_c_state[42];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[38];
  o_c_state[45] = i_c_state[28];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Back_counterclockwise;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[0];
  o_c_state[1] = i_c_state[1];
  o_c_state[2] = i_c_state[8];
  o_c_state[3] = i_c_state[23];
  o_c_state[4] = i_c_state[21];
  o_c_state[5] = i_c_state[5];
  o_c_state[6] = i_c_state[6];
  o_c_state[7] = i_c_state[4];
  o_c_state[8] = i_c_state[14];
  o_c_state[9] = i_c_state[9];
  o_c_state[10] = i_c_state[3];
  o_c_state[11] = i_c_state[11];
  o_c_state[12] = i_c_state[12];
  o_c_state[13] = i_c_state[10];
  o_c_state[14] = i_c_state[20];
  o_c_state[15] = i_c_state[15];
  o_c_state[16] = i_c_state[16];
  o_c_state[17] = i_c_state[7];
  o_c_state[18] = i_c_state[18];
  o_c_state[19] = i_c_state[19];
  o_c_state[20] = i_c_state[2];
  o_c_state[21] = i_c_state[17];
  o_c_state[22] = i_c_state[22];
  o_c_state[23] = i_c_state[13];
  o_c_state[24] = i_c_state[24];
  o_c_state[25] = i_c_state[25];
  o_c_state[26] = i_c_state[32];
  o_c_state[27] = i_c_state[27];
  o_c_state[28] = i_c_state[45];
  o_c_state[29] = i_c_state[29];
  o_c_state[30] = i_c_state[30];
  o_c_state[31] = i_c_state[28];
  o_c_state[32] = i_c_state[38];
  o_c_state[33] = i_c_state[33];
  o_c_state[34] = i_c_state[34];
  o_c_state[35] = i_c_state[35];
  o_c_state[36] = i_c_state[36];
  o_c_state[37] = i_c_state[37];
  o_c_state[38] = i_c_state[44];
  o_c_state[39] = i_c_state[39];
  o_c_state[40] = i_c_state[40];
  o_c_state[41] = i_c_state[31];
  o_c_state[42] = i_c_state[42];
  o_c_state[43] = i_c_state[43];
  o_c_state[44] = i_c_state[26];
  o_c_state[45] = i_c_state[41];
  o_c_state[46] = i_c_state[46];
  o_c_state[47] = i_c_state[47];
  end
  endtask
task Front_to_top;
  input [2:0] i_c_state [0:47];
 output [2:0] o_c_state[0:47];
 begin
  o_c_state[0] = i_c_state[5];
  o_c_state[1] = i_c_state[19];
  o_c_state[2] = i_c_state[16];
  o_c_state[3] = i_c_state[9];
  o_c_state[4] = i_c_state[0];
  o_c_state[5] = i_c_state[14];
  o_c_state[6] = i_c_state[11];
  o_c_state[7] = i_c_state[1];
  o_c_state[8] = i_c_state[22];
  o_c_state[9] = i_c_state[15];
  o_c_state[10] = i_c_state[6];
  o_c_state[11] = i_c_state[20];
  o_c_state[12] = i_c_state[17];
  o_c_state[13] = i_c_state[7];
  o_c_state[14] = i_c_state[4];
  o_c_state[15] = i_c_state[21];
  o_c_state[16] = i_c_state[12];
  o_c_state[17] = i_c_state[2];
  o_c_state[18] = i_c_state[23];
  o_c_state[19] = i_c_state[13];
  o_c_state[20] = i_c_state[10];
  o_c_state[21] = i_c_state[3];
  o_c_state[22] = i_c_state[18];
  o_c_state[23] = i_c_state[8];
  o_c_state[24] = i_c_state[29];
  o_c_state[25] = i_c_state[43];
  o_c_state[26] = i_c_state[40];
  o_c_state[27] = i_c_state[33];
  o_c_state[28] = i_c_state[24];
  o_c_state[29] = i_c_state[38];
  o_c_state[30] = i_c_state[35];
  o_c_state[31] = i_c_state[25];
  o_c_state[32] = i_c_state[46];
  o_c_state[33] = i_c_state[39];
  o_c_state[34] = i_c_state[30];
  o_c_state[35] = i_c_state[44];
  o_c_state[36] = i_c_state[41];
  o_c_state[37] = i_c_state[31];
  o_c_state[38] = i_c_state[28];
  o_c_state[39] = i_c_state[45];
  o_c_state[40] = i_c_state[36];
  o_c_state[41] = i_c_state[26];
  o_c_state[42] = i_c_state[47];
  o_c_state[43] = i_c_state[37];
  o_c_state[44] = i_c_state[34];
  o_c_state[45] = i_c_state[27];
  o_c_state[46] = i_c_state[42];
  o_c_state[47] = i_c_state[32];
  end
  endtask
